module iverilog_dump();
initial begin
    $dumpfile("tb_dllp_transmit.fst");
    $dumpvars(0, tb_dllp_transmit);
end
endmodule
