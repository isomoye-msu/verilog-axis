module block_alignment
  import pcie_phy_pkg::*;
#(
    // TLP data width
    parameter int DATA_WIDTH    = 32,
    // TLP strobe width
    // parameter int STRB_WIDTH    = DATA_WIDTH / 8,
    // parameter int KEEP_WIDTH    = STRB_WI1DTH,
    // parameter int USER_WIDTH    = 1,
    parameter int MAX_NUM_LANES = 4
) (
    //clocks and resets
    input  logic                                           clk_i,              // Clock signal
    input  logic                                           rst_i,              // Reset signal
    input  logic                                           phy_link_up_i,
    input  logic                                           lane_reverse_i,
    input  rate_speed_e                                    curr_data_rate_i,
    input  logic        [( MAX_NUM_LANES* DATA_WIDTH)-1:0] data_i,
    input  logic        [               MAX_NUM_LANES-1:0] data_valid_i,
    input  logic        [           (4*MAX_NUM_LANES)-1:0] data_k_i,
    input  logic        [           (2*MAX_NUM_LANES)-1:0] sync_header_i,
    output logic        [( MAX_NUM_LANES* DATA_WIDTH)-1:0] data_o,
    output logic        [               MAX_NUM_LANES-1:0] data_valid_o,
    output logic        [           (4*MAX_NUM_LANES)-1:0] data_k_o,
    output logic        [           (2*MAX_NUM_LANES)-1:0] sync_header_o,
    input  logic        [                             5:0] pipe_width_i,
    input  logic        [                             5:0] num_active_lanes_i
);



  localparam int PipeWidthGen1 = 8;
  localparam int PipeWidthGen2 = 16;
  localparam int PipeWidthGen3 = 16;
  localparam int PipeWidthGen4 = 32;
  localparam int PipeWidthGen5 = 32;
  localparam int BytesPerTransfer = DATA_WIDTH / 8;
  localparam int MaxWordsPerTransaction = 512 / DATA_WIDTH;

  // typedef enum logic [4:0] {
  //   ST_IDLE,
  //   ST_SEND_DATA,
  //   ST_LAST_DATA
  // } data_mux_st_e;


  // block_alignment_st_e                                    curr_state;
  // block_alignment_st_e                                    next_state;

  logic [( MAX_NUM_LANES* DATA_WIDTH)-1:0] data_c;
  logic [( MAX_NUM_LANES* DATA_WIDTH)-1:0] data_r;
  logic [               MAX_NUM_LANES-1:0] data_valid_c;
  logic [               MAX_NUM_LANES-1:0] data_valid_r;
  logic [           (4*MAX_NUM_LANES)-1:0] data_k_c;
  logic [           (4*MAX_NUM_LANES)-1:0] data_k_r;
  logic [           (2*MAX_NUM_LANES)-1:0] sync_header_c;
  logic [           (2*MAX_NUM_LANES)-1:0] sync_header_r;



  logic [                             5:0] word_count_c;
  logic [                             5:0] word_count_r;

  logic                                    is_ordered_set;
  logic                                    is_data;
  logic                                    ready_out;
  logic [                             7:0] lane_number;


  always_ff @(posedge clk_i) begin : main_seq_block
    if (rst_i) begin
      data_valid_r <= '0;
      // os_data_valid_r       <= '0;
      // tlp_dllp_data_valid_r <= '0;
    end else begin
      data_valid_r <= data_valid_c;
    end
    sync_header_r <= sync_header_c;
    data_k_r      <= data_k_c;
    data_r        <= data_c;
    // data_r                 <= data_c;
  end



  always_comb begin : block_alignment_combinational_logic
    data_c        = '0;
    data_valid_c  = '0;
    data_k_c      = '0;
    sync_header_c = '0;
    lane_number   = '0;
    if (phy_link_up_i) begin
      if (pipe_width_i == 8'd8 && |data_valid_i) begin
        for (int lane = 0; lane < MAX_NUM_LANES; lane++) begin
          lane_number = lane_reverse_i ? (num_active_lanes_i - 1) - lane : lane;
          if (lane < num_active_lanes_i) begin
            data_c[lane*8+:8] = data_i[BytesPerTransfer*lane_number*8+:8];
            data_valid_c[lane] = data_valid_i[lane_number];
            data_k_c[lane*4+:4] = data_k_i[BytesPerTransfer*lane_number*4+:4];
            sync_header_c[lane*2+:2] = sync_header_i[lane_number*2+:2];
          end
        end
      end
    end
  end


  assign sync_header_o = sync_header_r;
  assign data_valid_o  = data_valid_r;
  assign data_k_o      = data_k_r;
  assign data_o        = data_r;
endmodule
